library ieee;
use ieee.std_logic_1164.all;

use work.skinnypkg.all;

attribute S          : string;
attribute KEEP       : string;
attribute SYN_KEEP   : string;

entity g is
	port (x0, x1, x2, x3 : in  std_logic_vector(8 downto 0);
          y0, y1, y2, y3 : out std_logic_vector(7 downto 0));

    attribute S        of y0, y1, y2, y3  : signal is "true";
    attribute KEEP     of y0, y1, y2, y3  : signal is "true";
    attribute SYN_KEEP of y0, y1, y2, y3  : signal is "true";
end g;

attribute S        of g : entity is "true";
attribute KEEP     of g : entity is "true";
attribute SYN_KEEP of g : entity is "true";

architecture structural of g is
 
    signal w0, w1, w2, w3 : std_logic_vector(7 downto 0);

    attribute S        of w0, w1, w2, w3  : signal is "true";
    attribute KEEP     of w0, w1, w2, w3  : signal is "true";
    attribute SYN_KEEP of w0, w1, w2, w3  : signal is "true";

    attribute S        of p0, p1, p2, p3  : label is "true";
    attribute KEEP     of p0, p1, p2, p3  : label is "true";
    attribute SYN_KEEP of p0, p1, p2, p3  : label is "true";

begin

	p0 : entity work.g0 port map (
        x1(0), x2(0), x3(0),
        x1(1), x2(1), x3(1),
        x1(2), x2(2), x3(2),
        x1(3), x2(3), x3(3),
        x1(4), x2(4), x3(4),
        x1(5), x2(5), x3(5),
        x1(6), x2(6), x3(6),
        x1(7), x2(7), x3(7),
        x1(8), x2(8), x3(8),

        w0(0), w0(1), w0(2), w0(3), w0(4), w0(5), w0(6), w0(7)
    );
	
    p1 : entity work.g1 port map (
        x0(0), x2(0), x3(0),
        x0(1), x2(1), x3(1),
        x0(2), x2(2), x3(2),
        x0(3), x2(3), x3(3),
        x0(4), x2(4), x3(4),
        x0(5), x2(5), x3(5),
        x0(6), x2(6), x3(6),
        x0(7), x2(7), x3(7),
        x0(8), x2(8), x3(8),

        w1(0), w1(1), w1(2), w1(3), w1(4), w1(5), w1(6), w1(7)
    );
    
    p2 : entity work.g2 port map (
        x0(0), x1(0), x3(0),
        x0(1), x1(1), x3(1),
        x0(2), x1(2), x3(2),
        x0(3), x1(3), x3(3),
        x0(4), x1(4), x3(4),
        x0(5), x1(5), x3(5),
        x0(6), x1(6), x3(6),
        x0(7), x1(7), x3(7),
        x0(8), x1(8), x3(8),

        w2(0), w2(1), w2(2), w2(3), w2(4), w2(5), w2(6), w2(7)
    );
    
    p3 : entity work.g3 port map (
        x0(0), x1(0), x2(0),
        x0(1), x1(1), x2(1),
        x0(2), x1(2), x2(2),
        x0(3), x1(3), x2(3),
        x0(4), x1(4), x2(4),
        x0(5), x1(5), x2(5),
        x0(6), x1(6), x2(6),
        x0(7), x1(7), x2(7),
        x0(8), x1(8), x2(8),

        w3(0), w3(1), w3(2), w3(3), w3(4), w3(5), w3(6), w3(7)
    );
    
    y0 <= w0;
    y1 <= w1;
    y2 <= w2;
    y3 <= w3;

end structural;
